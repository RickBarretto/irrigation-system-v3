module select_led_color (
    // R, G, B
    output [2:0] color,

    input cleaning,
    input adubation,
    input error
);

endmodule