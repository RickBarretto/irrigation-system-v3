module tank_empting_decoder (
    output [6:0] column_4,
    output [6:0] column_3,
    output [6:0] column_2,
    output [6:0] column_1,
    output [6:0] column_0,

    // 3bits encoded counter
    input [2:0] water_level
);

endmodule