module tank_cleaning_decoder (
    output [6:0] column_2,
    output [6:0] column_1,
    output [6:0] column_0
);

endmodule